/*
 * bp_pce_pkg.vh
 *
 * This file contains the interface structures used for communication 
 * between BlackParrot and OpenPiton
 *
 */

package bp_pce_pkg;

  `include "bp_pce_l15_if.svh"

endpackage : bp_pce_pkg
